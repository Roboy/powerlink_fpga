// soc_system.v

// Generated using ACDS version 14.0 200 at 2017.06.23.23:56:49

`timescale 1 ps / 1 ps
module soc_system (
		input  wire        clk50_clk,                           //                  clk50.clk
		input  wire        clk100_clk,                          //                 clk100.clk
		input  wire [7:0]  node_switch_pio_export,              //        node_switch_pio.export
		input  wire        clk25_clk,                           //                  clk25.clk
		output wire [7:0]  pcp_0_benchmark_pio_export,          //    pcp_0_benchmark_pio.export
		input  wire        reset_reset_n,                       //                  reset.reset_n
		output wire [20:0] tri_state_0_tcm_address_out,         //            tri_state_0.tcm_address_out
		output wire [1:0]  tri_state_0_tcm_byteenable_n_out,    //                       .tcm_byteenable_n_out
		output wire [0:0]  tri_state_0_tcm_read_n_out,          //                       .tcm_read_n_out
		output wire [0:0]  tri_state_0_tcm_write_n_out,         //                       .tcm_write_n_out
		inout  wire [15:0] tri_state_0_tcm_data_out,            //                       .tcm_data_out
		output wire [0:0]  tri_state_0_tcm_chipselect_n_out,    //                       .tcm_chipselect_n_out
		output wire [1:0]  openmac_0_mii_txEnable,              //          openmac_0_mii.txEnable
		output wire [7:0]  openmac_0_mii_txData,                //                       .txData
		input  wire [1:0]  openmac_0_mii_txClk,                 //                       .txClk
		input  wire [1:0]  openmac_0_mii_rxError,               //                       .rxError
		input  wire [1:0]  openmac_0_mii_rxDataValid,           //                       .rxDataValid
		input  wire [7:0]  openmac_0_mii_rxData,                //                       .rxData
		input  wire [1:0]  openmac_0_mii_rxClk,                 //                       .rxClk
		output wire [1:0]  openmac_0_smi_nPhyRst,               //          openmac_0_smi.nPhyRst
		output wire [1:0]  openmac_0_smi_clk,                   //                       .clk
		inout  wire [1:0]  openmac_0_smi_dio,                   //                       .dio
		input  wire        pcp_0_cpu_resetrequest_resetrequest, // pcp_0_cpu_resetrequest.resetrequest
		output wire        pcp_0_cpu_resetrequest_resettaken,   //                       .resettaken
		output wire [1:0]  powerlink_led_export,                //          powerlink_led.export
		input  wire [31:0] app_pio_in_port,                     //                app_pio.in_port
		output wire [31:0] app_pio_out_port,                    //                       .out_port
		output wire        openmac_0_pktactivity_export         //  openmac_0_pktactivity.export
	);

	wire         sram_0_tcm_chipselect_n_out;                                          // sram_0:tcm_chipselect_n_out -> tri_state_0:tcs_tcm_chipselect_n_out
	wire         sram_0_tcm_grant;                                                     // tri_state_0:grant -> sram_0:tcm_grant
	wire         sram_0_tcm_data_outen;                                                // sram_0:tcm_data_outen -> tri_state_0:tcs_tcm_data_outen
	wire         sram_0_tcm_request;                                                   // sram_0:tcm_request -> tri_state_0:request
	wire  [15:0] sram_0_tcm_data_out;                                                  // sram_0:tcm_data_out -> tri_state_0:tcs_tcm_data_out
	wire         sram_0_tcm_write_n_out;                                               // sram_0:tcm_write_n_out -> tri_state_0:tcs_tcm_write_n_out
	wire  [20:0] sram_0_tcm_address_out;                                               // sram_0:tcm_address_out -> tri_state_0:tcs_tcm_address_out
	wire  [15:0] sram_0_tcm_data_in;                                                   // tri_state_0:tcs_tcm_data_in -> sram_0:tcm_data_in
	wire   [1:0] sram_0_tcm_byteenable_n_out;                                          // sram_0:tcm_byteenable_n_out -> tri_state_0:tcs_tcm_byteenable_n_out
	wire         sram_0_tcm_read_n_out;                                                // sram_0:tcm_read_n_out -> tri_state_0:tcs_tcm_read_n_out
	wire   [0:0] pcp_0_slow_bridge_burstcount;                                         // pcp_0:slow_bridge_burstcount -> mm_interconnect_0:pcp_0_slow_bridge_burstcount
	wire         pcp_0_slow_bridge_waitrequest;                                        // mm_interconnect_0:pcp_0_slow_bridge_waitrequest -> pcp_0:slow_bridge_waitrequest
	wire  [14:0] pcp_0_slow_bridge_address;                                            // pcp_0:slow_bridge_address -> mm_interconnect_0:pcp_0_slow_bridge_address
	wire  [31:0] pcp_0_slow_bridge_writedata;                                          // pcp_0:slow_bridge_writedata -> mm_interconnect_0:pcp_0_slow_bridge_writedata
	wire         pcp_0_slow_bridge_write;                                              // pcp_0:slow_bridge_write -> mm_interconnect_0:pcp_0_slow_bridge_write
	wire         pcp_0_slow_bridge_read;                                               // pcp_0:slow_bridge_read -> mm_interconnect_0:pcp_0_slow_bridge_read
	wire  [31:0] pcp_0_slow_bridge_readdata;                                           // mm_interconnect_0:pcp_0_slow_bridge_readdata -> pcp_0:slow_bridge_readdata
	wire         pcp_0_slow_bridge_debugaccess;                                        // pcp_0:slow_bridge_debugaccess -> mm_interconnect_0:pcp_0_slow_bridge_debugaccess
	wire   [3:0] pcp_0_slow_bridge_byteenable;                                         // pcp_0:slow_bridge_byteenable -> mm_interconnect_0:pcp_0_slow_bridge_byteenable
	wire         pcp_0_slow_bridge_readdatavalid;                                      // mm_interconnect_0:pcp_0_slow_bridge_readdatavalid -> pcp_0:slow_bridge_readdatavalid
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;                        // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;                       // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [1:0] mm_interconnect_0_node_switch_pio_s1_address;                         // mm_interconnect_0:node_switch_pio_s1_address -> node_switch_pio:address
	wire  [31:0] mm_interconnect_0_node_switch_pio_s1_readdata;                        // node_switch_pio:readdata -> mm_interconnect_0:node_switch_pio_s1_readdata
	wire         mm_interconnect_0_openmac_0_mactimer_waitrequest;                     // openmac_0:avs_macTimer_waitrequest -> mm_interconnect_0:openmac_0_macTimer_waitrequest
	wire  [31:0] mm_interconnect_0_openmac_0_mactimer_writedata;                       // mm_interconnect_0:openmac_0_macTimer_writedata -> openmac_0:avs_macTimer_writedata
	wire   [2:0] mm_interconnect_0_openmac_0_mactimer_address;                         // mm_interconnect_0:openmac_0_macTimer_address -> openmac_0:avs_macTimer_address
	wire         mm_interconnect_0_openmac_0_mactimer_chipselect;                      // mm_interconnect_0:openmac_0_macTimer_chipselect -> openmac_0:avs_macTimer_chipselect
	wire         mm_interconnect_0_openmac_0_mactimer_write;                           // mm_interconnect_0:openmac_0_macTimer_write -> openmac_0:avs_macTimer_write
	wire         mm_interconnect_0_openmac_0_mactimer_read;                            // mm_interconnect_0:openmac_0_macTimer_read -> openmac_0:avs_macTimer_read
	wire  [31:0] mm_interconnect_0_openmac_0_mactimer_readdata;                        // openmac_0:avs_macTimer_readdata -> mm_interconnect_0:openmac_0_macTimer_readdata
	wire   [3:0] mm_interconnect_0_openmac_0_mactimer_byteenable;                      // mm_interconnect_0:openmac_0_macTimer_byteenable -> openmac_0:avs_macTimer_byteenable
	wire         mm_interconnect_0_openmac_0_macreg_waitrequest;                       // openmac_0:avs_macReg_waitrequest -> mm_interconnect_0:openmac_0_macReg_waitrequest
	wire  [15:0] mm_interconnect_0_openmac_0_macreg_writedata;                         // mm_interconnect_0:openmac_0_macReg_writedata -> openmac_0:avs_macReg_writedata
	wire  [11:0] mm_interconnect_0_openmac_0_macreg_address;                           // mm_interconnect_0:openmac_0_macReg_address -> openmac_0:avs_macReg_address
	wire         mm_interconnect_0_openmac_0_macreg_chipselect;                        // mm_interconnect_0:openmac_0_macReg_chipselect -> openmac_0:avs_macReg_chipselect
	wire         mm_interconnect_0_openmac_0_macreg_write;                             // mm_interconnect_0:openmac_0_macReg_write -> openmac_0:avs_macReg_write
	wire         mm_interconnect_0_openmac_0_macreg_read;                              // mm_interconnect_0:openmac_0_macReg_read -> openmac_0:avs_macReg_read
	wire  [15:0] mm_interconnect_0_openmac_0_macreg_readdata;                          // openmac_0:avs_macReg_readdata -> mm_interconnect_0:openmac_0_macReg_readdata
	wire   [1:0] mm_interconnect_0_openmac_0_macreg_byteenable;                        // mm_interconnect_0:openmac_0_macReg_byteenable -> openmac_0:avs_macReg_byteenable
	wire  [31:0] mm_interconnect_0_app_pio_s1_writedata;                               // mm_interconnect_0:app_pio_s1_writedata -> app_pio:writedata
	wire   [1:0] mm_interconnect_0_app_pio_s1_address;                                 // mm_interconnect_0:app_pio_s1_address -> app_pio:address
	wire         mm_interconnect_0_app_pio_s1_chipselect;                              // mm_interconnect_0:app_pio_s1_chipselect -> app_pio:chipselect
	wire         mm_interconnect_0_app_pio_s1_write;                                   // mm_interconnect_0:app_pio_s1_write -> app_pio:write_n
	wire  [31:0] mm_interconnect_0_app_pio_s1_readdata;                                // app_pio:readdata -> mm_interconnect_0:app_pio_s1_readdata
	wire   [0:0] pcp_0_cpu_bridge_burstcount;                                          // pcp_0:cpu_bridge_burstcount -> mm_interconnect_1:pcp_0_cpu_bridge_burstcount
	wire         pcp_0_cpu_bridge_waitrequest;                                         // mm_interconnect_1:pcp_0_cpu_bridge_waitrequest -> pcp_0:cpu_bridge_waitrequest
	wire  [21:0] pcp_0_cpu_bridge_address;                                             // pcp_0:cpu_bridge_address -> mm_interconnect_1:pcp_0_cpu_bridge_address
	wire  [31:0] pcp_0_cpu_bridge_writedata;                                           // pcp_0:cpu_bridge_writedata -> mm_interconnect_1:pcp_0_cpu_bridge_writedata
	wire         pcp_0_cpu_bridge_write;                                               // pcp_0:cpu_bridge_write -> mm_interconnect_1:pcp_0_cpu_bridge_write
	wire         pcp_0_cpu_bridge_read;                                                // pcp_0:cpu_bridge_read -> mm_interconnect_1:pcp_0_cpu_bridge_read
	wire  [31:0] pcp_0_cpu_bridge_readdata;                                            // mm_interconnect_1:pcp_0_cpu_bridge_readdata -> pcp_0:cpu_bridge_readdata
	wire         pcp_0_cpu_bridge_debugaccess;                                         // pcp_0:cpu_bridge_debugaccess -> mm_interconnect_1:pcp_0_cpu_bridge_debugaccess
	wire   [3:0] pcp_0_cpu_bridge_byteenable;                                          // pcp_0:cpu_bridge_byteenable -> mm_interconnect_1:pcp_0_cpu_bridge_byteenable
	wire         pcp_0_cpu_bridge_readdatavalid;                                       // mm_interconnect_1:pcp_0_cpu_bridge_readdatavalid -> pcp_0:cpu_bridge_readdatavalid
	wire  [13:0] openmac_0_dma_burstcount;                                             // openmac_0:avm_dma_burstcount -> mm_interconnect_1:openmac_0_dma_burstcount
	wire         openmac_0_dma_waitrequest;                                            // mm_interconnect_1:openmac_0_dma_waitrequest -> openmac_0:avm_dma_waitrequest
	wire  [15:0] openmac_0_dma_writedata;                                              // openmac_0:avm_dma_writedata -> mm_interconnect_1:openmac_0_dma_writedata
	wire  [20:0] openmac_0_dma_address;                                                // openmac_0:avm_dma_address -> mm_interconnect_1:openmac_0_dma_address
	wire         openmac_0_dma_write;                                                  // openmac_0:avm_dma_write -> mm_interconnect_1:openmac_0_dma_write
	wire         openmac_0_dma_read;                                                   // openmac_0:avm_dma_read -> mm_interconnect_1:openmac_0_dma_read
	wire  [15:0] openmac_0_dma_readdata;                                               // mm_interconnect_1:openmac_0_dma_readdata -> openmac_0:avm_dma_readdata
	wire   [1:0] openmac_0_dma_byteenable;                                             // openmac_0:avm_dma_byteenable -> mm_interconnect_1:openmac_0_dma_byteenable
	wire         openmac_0_dma_readdatavalid;                                          // mm_interconnect_1:openmac_0_dma_readdatavalid -> openmac_0:avm_dma_readdatavalid
	wire         mm_interconnect_1_sram_0_uas_waitrequest;                             // sram_0:uas_waitrequest -> mm_interconnect_1:sram_0_uas_waitrequest
	wire   [1:0] mm_interconnect_1_sram_0_uas_burstcount;                              // mm_interconnect_1:sram_0_uas_burstcount -> sram_0:uas_burstcount
	wire  [15:0] mm_interconnect_1_sram_0_uas_writedata;                               // mm_interconnect_1:sram_0_uas_writedata -> sram_0:uas_writedata
	wire  [20:0] mm_interconnect_1_sram_0_uas_address;                                 // mm_interconnect_1:sram_0_uas_address -> sram_0:uas_address
	wire         mm_interconnect_1_sram_0_uas_lock;                                    // mm_interconnect_1:sram_0_uas_lock -> sram_0:uas_lock
	wire         mm_interconnect_1_sram_0_uas_write;                                   // mm_interconnect_1:sram_0_uas_write -> sram_0:uas_write
	wire         mm_interconnect_1_sram_0_uas_read;                                    // mm_interconnect_1:sram_0_uas_read -> sram_0:uas_read
	wire  [15:0] mm_interconnect_1_sram_0_uas_readdata;                                // sram_0:uas_readdata -> mm_interconnect_1:sram_0_uas_readdata
	wire         mm_interconnect_1_sram_0_uas_debugaccess;                             // mm_interconnect_1:sram_0_uas_debugaccess -> sram_0:uas_debugaccess
	wire         mm_interconnect_1_sram_0_uas_readdatavalid;                           // sram_0:uas_readdatavalid -> mm_interconnect_1:sram_0_uas_readdatavalid
	wire   [1:0] mm_interconnect_1_sram_0_uas_byteenable;                              // mm_interconnect_1:sram_0_uas_byteenable -> sram_0:uas_byteenable
	wire   [0:0] pcp_0_flash_bridge_burstcount;                                        // pcp_0:flash_bridge_burstcount -> mm_interconnect_2:pcp_0_flash_bridge_burstcount
	wire         pcp_0_flash_bridge_waitrequest;                                       // mm_interconnect_2:pcp_0_flash_bridge_waitrequest -> pcp_0:flash_bridge_waitrequest
	wire  [21:0] pcp_0_flash_bridge_address;                                           // pcp_0:flash_bridge_address -> mm_interconnect_2:pcp_0_flash_bridge_address
	wire  [31:0] pcp_0_flash_bridge_writedata;                                         // pcp_0:flash_bridge_writedata -> mm_interconnect_2:pcp_0_flash_bridge_writedata
	wire         pcp_0_flash_bridge_write;                                             // pcp_0:flash_bridge_write -> mm_interconnect_2:pcp_0_flash_bridge_write
	wire         pcp_0_flash_bridge_read;                                              // pcp_0:flash_bridge_read -> mm_interconnect_2:pcp_0_flash_bridge_read
	wire  [31:0] pcp_0_flash_bridge_readdata;                                          // mm_interconnect_2:pcp_0_flash_bridge_readdata -> pcp_0:flash_bridge_readdata
	wire         pcp_0_flash_bridge_debugaccess;                                       // pcp_0:flash_bridge_debugaccess -> mm_interconnect_2:pcp_0_flash_bridge_debugaccess
	wire   [3:0] pcp_0_flash_bridge_byteenable;                                        // pcp_0:flash_bridge_byteenable -> mm_interconnect_2:pcp_0_flash_bridge_byteenable
	wire         pcp_0_flash_bridge_readdatavalid;                                     // mm_interconnect_2:pcp_0_flash_bridge_readdatavalid -> pcp_0:flash_bridge_readdatavalid
	wire  [31:0] mm_interconnect_2_epcs_flash_controller_epcs_control_port_writedata;  // mm_interconnect_2:epcs_flash_controller_epcs_control_port_writedata -> epcs_flash_controller:writedata
	wire   [8:0] mm_interconnect_2_epcs_flash_controller_epcs_control_port_address;    // mm_interconnect_2:epcs_flash_controller_epcs_control_port_address -> epcs_flash_controller:address
	wire         mm_interconnect_2_epcs_flash_controller_epcs_control_port_chipselect; // mm_interconnect_2:epcs_flash_controller_epcs_control_port_chipselect -> epcs_flash_controller:chipselect
	wire         mm_interconnect_2_epcs_flash_controller_epcs_control_port_write;      // mm_interconnect_2:epcs_flash_controller_epcs_control_port_write -> epcs_flash_controller:write_n
	wire         mm_interconnect_2_epcs_flash_controller_epcs_control_port_read;       // mm_interconnect_2:epcs_flash_controller_epcs_control_port_read -> epcs_flash_controller:read_n
	wire  [31:0] mm_interconnect_2_epcs_flash_controller_epcs_control_port_readdata;   // epcs_flash_controller:readdata -> mm_interconnect_2:epcs_flash_controller_epcs_control_port_readdata
	wire         irq_mapper_receiver0_irq;                                             // openmac_0:ins_timerIrq_irq -> irq_mapper:receiver0_irq
	wire   [0:0] pcp_0_sync_irq_irq;                                                   // irq_mapper:sender_irq -> pcp_0:sync_irq_irq
	wire         irq_mapper_001_receiver0_irq;                                         // openmac_0:ins_macIrq_irq -> irq_mapper_001:receiver0_irq
	wire   [0:0] pcp_0_mac_irq_irq;                                                    // irq_mapper_001:sender_irq -> pcp_0:mac_irq_irq
	wire         irq_mapper_002_receiver0_irq;                                         // epcs_flash_controller:irq -> irq_mapper_002:receiver0_irq
	wire   [3:0] pcp_0_gp_irq_irq;                                                     // irq_mapper_002:sender_irq -> pcp_0:gp_irq_irq
	wire         rst_controller_reset_out_reset;                                       // rst_controller:reset_out -> [app_pio:reset_n, irq_mapper:reset, irq_mapper_001:reset, irq_mapper_002:reset, mm_interconnect_0:pcp_0_rst_clk50_reset_bridge_in_reset_reset, mm_interconnect_0:sysid_reset_reset_bridge_in_reset_reset, mm_interconnect_2:pcp_0_flash_bridge_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_2:pcp_0_rst_clk50_reset_bridge_in_reset_reset, node_switch_pio:reset_n, sysid:reset_n]
	wire         rst_controller_001_reset_out_reset;                                   // rst_controller_001:reset_out -> pcp_0:rst_clk50_reset_n
	wire         rst_controller_002_reset_out_reset;                                   // rst_controller_002:reset_out -> pcp_0:rst_clk100_reset_n
	wire         rst_controller_003_reset_out_reset;                                   // rst_controller_003:reset_out -> [mm_interconnect_1:pcp_0_rst_clk50_reset_bridge_in_reset_reset, mm_interconnect_1:sram_0_reset_reset_bridge_in_reset_reset, sram_0:reset_reset, tri_state_0:reset]
	wire         rst_controller_004_reset_out_reset;                                   // rst_controller_004:reset_out -> openmac_0:rsi_mainRst_reset
	wire         rst_controller_005_reset_out_reset;                                   // rst_controller_005:reset_out -> openmac_0:rsi_dmaRst_reset
	wire         rst_controller_006_reset_out_reset;                                   // rst_controller_006:reset_out -> [epcs_flash_controller:reset_n, mm_interconnect_2:epcs_flash_controller_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_006_reset_out_reset_req;                               // rst_controller_006:reset_req -> epcs_flash_controller:reset_req
	wire         pcp_0_jtag_reset_reset;                                               // pcp_0:jtag_reset_reset -> rst_controller_006:reset_in3

	soc_system_node_switch_pio node_switch_pio (
		.clk      (clk50_clk),                                     //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_0_node_switch_pio_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_node_switch_pio_s1_readdata), //                    .readdata
		.in_port  (node_switch_pio_export)                         // external_connection.export
	);

	soc_system_pcp_0 pcp_0 (
		.clk50_clk                     (clk50_clk),                           //            clk50.clk
		.rst_clk50_reset_n             (~rst_controller_001_reset_out_reset), //        rst_clk50.reset_n
		.clk100_clk                    (clk100_clk),                          //           clk100.clk
		.rst_clk100_reset_n            (~rst_controller_002_reset_out_reset), //       rst_clk100.reset_n
		.benchmark_pio_export          (pcp_0_benchmark_pio_export),          //    benchmark_pio.export
		.cpu_bridge_waitrequest        (pcp_0_cpu_bridge_waitrequest),        //       cpu_bridge.waitrequest
		.cpu_bridge_readdata           (pcp_0_cpu_bridge_readdata),           //                 .readdata
		.cpu_bridge_readdatavalid      (pcp_0_cpu_bridge_readdatavalid),      //                 .readdatavalid
		.cpu_bridge_burstcount         (pcp_0_cpu_bridge_burstcount),         //                 .burstcount
		.cpu_bridge_writedata          (pcp_0_cpu_bridge_writedata),          //                 .writedata
		.cpu_bridge_address            (pcp_0_cpu_bridge_address),            //                 .address
		.cpu_bridge_write              (pcp_0_cpu_bridge_write),              //                 .write
		.cpu_bridge_read               (pcp_0_cpu_bridge_read),               //                 .read
		.cpu_bridge_byteenable         (pcp_0_cpu_bridge_byteenable),         //                 .byteenable
		.cpu_bridge_debugaccess        (pcp_0_cpu_bridge_debugaccess),        //                 .debugaccess
		.slow_bridge_waitrequest       (pcp_0_slow_bridge_waitrequest),       //      slow_bridge.waitrequest
		.slow_bridge_readdata          (pcp_0_slow_bridge_readdata),          //                 .readdata
		.slow_bridge_readdatavalid     (pcp_0_slow_bridge_readdatavalid),     //                 .readdatavalid
		.slow_bridge_burstcount        (pcp_0_slow_bridge_burstcount),        //                 .burstcount
		.slow_bridge_writedata         (pcp_0_slow_bridge_writedata),         //                 .writedata
		.slow_bridge_address           (pcp_0_slow_bridge_address),           //                 .address
		.slow_bridge_write             (pcp_0_slow_bridge_write),             //                 .write
		.slow_bridge_read              (pcp_0_slow_bridge_read),              //                 .read
		.slow_bridge_byteenable        (pcp_0_slow_bridge_byteenable),        //                 .byteenable
		.slow_bridge_debugaccess       (pcp_0_slow_bridge_debugaccess),       //                 .debugaccess
		.sync_irq_irq                  (pcp_0_sync_irq_irq),                  //         sync_irq.irq
		.mac_irq_irq                   (pcp_0_mac_irq_irq),                   //          mac_irq.irq
		.flash_bridge_waitrequest      (pcp_0_flash_bridge_waitrequest),      //     flash_bridge.waitrequest
		.flash_bridge_readdata         (pcp_0_flash_bridge_readdata),         //                 .readdata
		.flash_bridge_readdatavalid    (pcp_0_flash_bridge_readdatavalid),    //                 .readdatavalid
		.flash_bridge_burstcount       (pcp_0_flash_bridge_burstcount),       //                 .burstcount
		.flash_bridge_writedata        (pcp_0_flash_bridge_writedata),        //                 .writedata
		.flash_bridge_address          (pcp_0_flash_bridge_address),          //                 .address
		.flash_bridge_write            (pcp_0_flash_bridge_write),            //                 .write
		.flash_bridge_read             (pcp_0_flash_bridge_read),             //                 .read
		.flash_bridge_byteenable       (pcp_0_flash_bridge_byteenable),       //                 .byteenable
		.flash_bridge_debugaccess      (pcp_0_flash_bridge_debugaccess),      //                 .debugaccess
		.gp_irq_irq                    (pcp_0_gp_irq_irq),                    //           gp_irq.irq
		.cpu_resetrequest_resetrequest (pcp_0_cpu_resetrequest_resetrequest), // cpu_resetrequest.resetrequest
		.cpu_resetrequest_resettaken   (pcp_0_cpu_resetrequest_resettaken),   //                 .resettaken
		.jtag_reset_reset              (pcp_0_jtag_reset_reset),              //       jtag_reset.reset
		.powerlink_led_export          (powerlink_led_export)                 //    powerlink_led.export
	);

	soc_system_sysid sysid (
		.clock    (clk50_clk),                                      //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	soc_system_sram_0 #(
		.TCM_ADDRESS_W                  (21),
		.TCM_DATA_W                     (16),
		.TCM_BYTEENABLE_W               (2),
		.TCM_READ_WAIT                  (1),
		.TCM_WRITE_WAIT                 (0),
		.TCM_SETUP_WAIT                 (0),
		.TCM_DATA_HOLD                  (0),
		.TCM_TURNAROUND_TIME            (1),
		.TCM_TIMING_UNITS               (1),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (2),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (1),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (1),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (0),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (1),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (1),
		.ACTIVE_LOW_OUTPUTENABLE        (0),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (0)
	) sram_0 (
		.clk_clk              (clk100_clk),                                 //   clk.clk
		.reset_reset          (rst_controller_003_reset_out_reset),         // reset.reset
		.uas_address          (mm_interconnect_1_sram_0_uas_address),       //   uas.address
		.uas_burstcount       (mm_interconnect_1_sram_0_uas_burstcount),    //      .burstcount
		.uas_read             (mm_interconnect_1_sram_0_uas_read),          //      .read
		.uas_write            (mm_interconnect_1_sram_0_uas_write),         //      .write
		.uas_waitrequest      (mm_interconnect_1_sram_0_uas_waitrequest),   //      .waitrequest
		.uas_readdatavalid    (mm_interconnect_1_sram_0_uas_readdatavalid), //      .readdatavalid
		.uas_byteenable       (mm_interconnect_1_sram_0_uas_byteenable),    //      .byteenable
		.uas_readdata         (mm_interconnect_1_sram_0_uas_readdata),      //      .readdata
		.uas_writedata        (mm_interconnect_1_sram_0_uas_writedata),     //      .writedata
		.uas_lock             (mm_interconnect_1_sram_0_uas_lock),          //      .lock
		.uas_debugaccess      (mm_interconnect_1_sram_0_uas_debugaccess),   //      .debugaccess
		.tcm_write_n_out      (sram_0_tcm_write_n_out),                     //   tcm.write_n_out
		.tcm_read_n_out       (sram_0_tcm_read_n_out),                      //      .read_n_out
		.tcm_chipselect_n_out (sram_0_tcm_chipselect_n_out),                //      .chipselect_n_out
		.tcm_request          (sram_0_tcm_request),                         //      .request
		.tcm_grant            (sram_0_tcm_grant),                           //      .grant
		.tcm_address_out      (sram_0_tcm_address_out),                     //      .address_out
		.tcm_byteenable_n_out (sram_0_tcm_byteenable_n_out),                //      .byteenable_n_out
		.tcm_data_out         (sram_0_tcm_data_out),                        //      .data_out
		.tcm_data_outen       (sram_0_tcm_data_outen),                      //      .data_outen
		.tcm_data_in          (sram_0_tcm_data_in)                          //      .data_in
	);

	soc_system_tri_state_0 tri_state_0 (
		.clk                      (clk100_clk),                         //   clk.clk
		.reset                    (rst_controller_003_reset_out_reset), // reset.reset
		.request                  (sram_0_tcm_request),                 //   tcs.request
		.grant                    (sram_0_tcm_grant),                   //      .grant
		.tcs_tcm_address_out      (sram_0_tcm_address_out),             //      .address_out
		.tcs_tcm_byteenable_n_out (sram_0_tcm_byteenable_n_out),        //      .byteenable_n_out
		.tcs_tcm_read_n_out       (sram_0_tcm_read_n_out),              //      .read_n_out
		.tcs_tcm_write_n_out      (sram_0_tcm_write_n_out),             //      .write_n_out
		.tcs_tcm_data_out         (sram_0_tcm_data_out),                //      .data_out
		.tcs_tcm_data_outen       (sram_0_tcm_data_outen),              //      .data_outen
		.tcs_tcm_data_in          (sram_0_tcm_data_in),                 //      .data_in
		.tcs_tcm_chipselect_n_out (sram_0_tcm_chipselect_n_out),        //      .chipselect_n_out
		.tcm_address_out          (tri_state_0_tcm_address_out),        //   out.tcm_address_out
		.tcm_byteenable_n_out     (tri_state_0_tcm_byteenable_n_out),   //      .tcm_byteenable_n_out
		.tcm_read_n_out           (tri_state_0_tcm_read_n_out),         //      .tcm_read_n_out
		.tcm_write_n_out          (tri_state_0_tcm_write_n_out),        //      .tcm_write_n_out
		.tcm_data_out             (tri_state_0_tcm_data_out),           //      .tcm_data_out
		.tcm_chipselect_n_out     (tri_state_0_tcm_chipselect_n_out)    //      .tcm_chipselect_n_out
	);

	alteraOpenmacTop #(
		.gPhyPortCount          (2),
		.gPhyPortType           (2),
		.gSmiPortCount          (2),
		.gEndianness            ("little"),
		.gEnableActivity        (1),
		.gEnableDmaObserver     (1),
		.gDmaAddrWidth          (21),
		.gDmaDataWidth          (16),
		.gDmaBurstCountWidth    (14),
		.gDmaWriteBurstLength   (1),
		.gDmaReadBurstLength    (8),
		.gDmaWriteFifoLength    (16),
		.gDmaReadFifoLength     (16),
		.gPacketBufferLocTx     (2),
		.gPacketBufferLocRx     (2),
		.gPacketBufferLog2Size  (4),
		.gTimerEnablePulse      (0),
		.gTimerEnablePulseWidth (0),
		.gTimerPulseRegWidth    (10)
	) openmac_0 (
		.csi_mainClk_clock        (clk50_clk),                                        //     mainClk.clk
		.csi_mainClkx2_clock      (clk100_clk),                                       //   mainClkx2.clk
		.csi_dmaClk_clock         (clk100_clk),                                       //      dmaClk.clk
		.rsi_mainRst_reset        (rst_controller_004_reset_out_reset),               //     mainRst.reset
		.rsi_dmaRst_reset         (rst_controller_005_reset_out_reset),               //      dmaRst.reset
		.avs_macReg_chipselect    (mm_interconnect_0_openmac_0_macreg_chipselect),    //      macReg.chipselect
		.avs_macReg_write         (mm_interconnect_0_openmac_0_macreg_write),         //            .write
		.avs_macReg_read          (mm_interconnect_0_openmac_0_macreg_read),          //            .read
		.avs_macReg_waitrequest   (mm_interconnect_0_openmac_0_macreg_waitrequest),   //            .waitrequest
		.avs_macReg_byteenable    (mm_interconnect_0_openmac_0_macreg_byteenable),    //            .byteenable
		.avs_macReg_address       (mm_interconnect_0_openmac_0_macreg_address),       //            .address
		.avs_macReg_writedata     (mm_interconnect_0_openmac_0_macreg_writedata),     //            .writedata
		.avs_macReg_readdata      (mm_interconnect_0_openmac_0_macreg_readdata),      //            .readdata
		.avs_macTimer_chipselect  (mm_interconnect_0_openmac_0_mactimer_chipselect),  //    macTimer.chipselect
		.avs_macTimer_write       (mm_interconnect_0_openmac_0_mactimer_write),       //            .write
		.avs_macTimer_read        (mm_interconnect_0_openmac_0_mactimer_read),        //            .read
		.avs_macTimer_waitrequest (mm_interconnect_0_openmac_0_mactimer_waitrequest), //            .waitrequest
		.avs_macTimer_address     (mm_interconnect_0_openmac_0_mactimer_address),     //            .address
		.avs_macTimer_byteenable  (mm_interconnect_0_openmac_0_mactimer_byteenable),  //            .byteenable
		.avs_macTimer_writedata   (mm_interconnect_0_openmac_0_mactimer_writedata),   //            .writedata
		.avs_macTimer_readdata    (mm_interconnect_0_openmac_0_mactimer_readdata),    //            .readdata
		.avm_dma_write            (openmac_0_dma_write),                              //         dma.write
		.avm_dma_read             (openmac_0_dma_read),                               //            .read
		.avm_dma_waitrequest      (openmac_0_dma_waitrequest),                        //            .waitrequest
		.avm_dma_readdatavalid    (openmac_0_dma_readdatavalid),                      //            .readdatavalid
		.avm_dma_byteenable       (openmac_0_dma_byteenable),                         //            .byteenable
		.avm_dma_address          (openmac_0_dma_address),                            //            .address
		.avm_dma_burstcount       (openmac_0_dma_burstcount),                         //            .burstcount
		.avm_dma_writedata        (openmac_0_dma_writedata),                          //            .writedata
		.avm_dma_readdata         (openmac_0_dma_readdata),                           //            .readdata
		.ins_timerIrq_irq         (irq_mapper_receiver0_irq),                         //    timerIrq.irq
		.ins_macIrq_irq           (irq_mapper_001_receiver0_irq),                     //      macIrq.irq
		.coe_mii_txEnable         (openmac_0_mii_txEnable),                           //         mii.export
		.coe_mii_txData           (openmac_0_mii_txData),                             //            .export
		.coe_mii_txClk            (openmac_0_mii_txClk),                              //            .export
		.coe_mii_rxError          (openmac_0_mii_rxError),                            //            .export
		.coe_mii_rxDataValid      (openmac_0_mii_rxDataValid),                        //            .export
		.coe_mii_rxData           (openmac_0_mii_rxData),                             //            .export
		.coe_mii_rxClk            (openmac_0_mii_rxClk),                              //            .export
		.coe_smi_nPhyRst          (openmac_0_smi_nPhyRst),                            //         smi.export
		.coe_smi_clk              (openmac_0_smi_clk),                                //            .export
		.coe_smi_dio              (openmac_0_smi_dio),                                //            .export
		.coe_pktActivity          (openmac_0_pktactivity_export),                     // pktActivity.export
		.csi_pktClk_clock         (1'b0),                                             // (terminated)
		.rsi_pktRst_reset         (1'b0),                                             // (terminated)
		.avs_pktBuf_chipselect    (1'b0),                                             // (terminated)
		.avs_pktBuf_write         (1'b0),                                             // (terminated)
		.avs_pktBuf_read          (1'b0),                                             // (terminated)
		.avs_pktBuf_waitrequest   (),                                                 // (terminated)
		.avs_pktBuf_byteenable    (4'b0000),                                          // (terminated)
		.avs_pktBuf_address       (2'b00),                                            // (terminated)
		.avs_pktBuf_writedata     (32'b00000000000000000000000000000000),             // (terminated)
		.avs_pktBuf_readdata      (),                                                 // (terminated)
		.ins_timerPulse_irq       (),                                                 // (terminated)
		.coe_rmii_txEnable        (),                                                 // (terminated)
		.coe_rmii_txData          (),                                                 // (terminated)
		.coe_rmii_rxError         (2'b00),                                            // (terminated)
		.coe_rmii_rxCrsDataValid  (2'b00),                                            // (terminated)
		.coe_rmii_rxData          (4'b0000)                                           // (terminated)
	);

	soc_system_epcs_flash_controller epcs_flash_controller (
		.clk           (clk50_clk),                                                            //               clk.clk
		.reset_n       (~rst_controller_006_reset_out_reset),                                  //             reset.reset_n
		.reset_req     (rst_controller_006_reset_out_reset_req),                               //                  .reset_req
		.address       (mm_interconnect_2_epcs_flash_controller_epcs_control_port_address),    // epcs_control_port.address
		.chipselect    (mm_interconnect_2_epcs_flash_controller_epcs_control_port_chipselect), //                  .chipselect
		.dataavailable (),                                                                     //                  .dataavailable
		.endofpacket   (),                                                                     //                  .endofpacket
		.read_n        (~mm_interconnect_2_epcs_flash_controller_epcs_control_port_read),      //                  .read_n
		.readdata      (mm_interconnect_2_epcs_flash_controller_epcs_control_port_readdata),   //                  .readdata
		.readyfordata  (),                                                                     //                  .readyfordata
		.write_n       (~mm_interconnect_2_epcs_flash_controller_epcs_control_port_write),     //                  .write_n
		.writedata     (mm_interconnect_2_epcs_flash_controller_epcs_control_port_writedata),  //                  .writedata
		.irq           (irq_mapper_002_receiver0_irq)                                          //               irq.irq
	);

	soc_system_app_pio app_pio (
		.clk        (clk50_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_app_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_app_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_app_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_app_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_app_pio_s1_readdata),   //                    .readdata
		.in_port    (app_pio_in_port),                         // external_connection.export
		.out_port   (app_pio_out_port)                         //                    .export
	);

	soc_system_mm_interconnect_0 mm_interconnect_0 (
		.clk50_clk_clk                               (clk50_clk),                                        //                             clk50_clk.clk
		.pcp_0_rst_clk50_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                   // pcp_0_rst_clk50_reset_bridge_in_reset.reset
		.sysid_reset_reset_bridge_in_reset_reset     (rst_controller_reset_out_reset),                   //     sysid_reset_reset_bridge_in_reset.reset
		.pcp_0_slow_bridge_address                   (pcp_0_slow_bridge_address),                        //                     pcp_0_slow_bridge.address
		.pcp_0_slow_bridge_waitrequest               (pcp_0_slow_bridge_waitrequest),                    //                                      .waitrequest
		.pcp_0_slow_bridge_burstcount                (pcp_0_slow_bridge_burstcount),                     //                                      .burstcount
		.pcp_0_slow_bridge_byteenable                (pcp_0_slow_bridge_byteenable),                     //                                      .byteenable
		.pcp_0_slow_bridge_read                      (pcp_0_slow_bridge_read),                           //                                      .read
		.pcp_0_slow_bridge_readdata                  (pcp_0_slow_bridge_readdata),                       //                                      .readdata
		.pcp_0_slow_bridge_readdatavalid             (pcp_0_slow_bridge_readdatavalid),                  //                                      .readdatavalid
		.pcp_0_slow_bridge_write                     (pcp_0_slow_bridge_write),                          //                                      .write
		.pcp_0_slow_bridge_writedata                 (pcp_0_slow_bridge_writedata),                      //                                      .writedata
		.pcp_0_slow_bridge_debugaccess               (pcp_0_slow_bridge_debugaccess),                    //                                      .debugaccess
		.app_pio_s1_address                          (mm_interconnect_0_app_pio_s1_address),             //                            app_pio_s1.address
		.app_pio_s1_write                            (mm_interconnect_0_app_pio_s1_write),               //                                      .write
		.app_pio_s1_readdata                         (mm_interconnect_0_app_pio_s1_readdata),            //                                      .readdata
		.app_pio_s1_writedata                        (mm_interconnect_0_app_pio_s1_writedata),           //                                      .writedata
		.app_pio_s1_chipselect                       (mm_interconnect_0_app_pio_s1_chipselect),          //                                      .chipselect
		.node_switch_pio_s1_address                  (mm_interconnect_0_node_switch_pio_s1_address),     //                    node_switch_pio_s1.address
		.node_switch_pio_s1_readdata                 (mm_interconnect_0_node_switch_pio_s1_readdata),    //                                      .readdata
		.openmac_0_macReg_address                    (mm_interconnect_0_openmac_0_macreg_address),       //                      openmac_0_macReg.address
		.openmac_0_macReg_write                      (mm_interconnect_0_openmac_0_macreg_write),         //                                      .write
		.openmac_0_macReg_read                       (mm_interconnect_0_openmac_0_macreg_read),          //                                      .read
		.openmac_0_macReg_readdata                   (mm_interconnect_0_openmac_0_macreg_readdata),      //                                      .readdata
		.openmac_0_macReg_writedata                  (mm_interconnect_0_openmac_0_macreg_writedata),     //                                      .writedata
		.openmac_0_macReg_byteenable                 (mm_interconnect_0_openmac_0_macreg_byteenable),    //                                      .byteenable
		.openmac_0_macReg_waitrequest                (mm_interconnect_0_openmac_0_macreg_waitrequest),   //                                      .waitrequest
		.openmac_0_macReg_chipselect                 (mm_interconnect_0_openmac_0_macreg_chipselect),    //                                      .chipselect
		.openmac_0_macTimer_address                  (mm_interconnect_0_openmac_0_mactimer_address),     //                    openmac_0_macTimer.address
		.openmac_0_macTimer_write                    (mm_interconnect_0_openmac_0_mactimer_write),       //                                      .write
		.openmac_0_macTimer_read                     (mm_interconnect_0_openmac_0_mactimer_read),        //                                      .read
		.openmac_0_macTimer_readdata                 (mm_interconnect_0_openmac_0_mactimer_readdata),    //                                      .readdata
		.openmac_0_macTimer_writedata                (mm_interconnect_0_openmac_0_mactimer_writedata),   //                                      .writedata
		.openmac_0_macTimer_byteenable               (mm_interconnect_0_openmac_0_mactimer_byteenable),  //                                      .byteenable
		.openmac_0_macTimer_waitrequest              (mm_interconnect_0_openmac_0_mactimer_waitrequest), //                                      .waitrequest
		.openmac_0_macTimer_chipselect               (mm_interconnect_0_openmac_0_mactimer_chipselect),  //                                      .chipselect
		.sysid_control_slave_address                 (mm_interconnect_0_sysid_control_slave_address),    //                   sysid_control_slave.address
		.sysid_control_slave_readdata                (mm_interconnect_0_sysid_control_slave_readdata)    //                                      .readdata
	);

	soc_system_mm_interconnect_1 mm_interconnect_1 (
		.clk100_clk_clk                              (clk100_clk),                                 //                            clk100_clk.clk
		.pcp_0_rst_clk50_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),         // pcp_0_rst_clk50_reset_bridge_in_reset.reset
		.sram_0_reset_reset_bridge_in_reset_reset    (rst_controller_003_reset_out_reset),         //    sram_0_reset_reset_bridge_in_reset.reset
		.openmac_0_dma_address                       (openmac_0_dma_address),                      //                         openmac_0_dma.address
		.openmac_0_dma_waitrequest                   (openmac_0_dma_waitrequest),                  //                                      .waitrequest
		.openmac_0_dma_burstcount                    (openmac_0_dma_burstcount),                   //                                      .burstcount
		.openmac_0_dma_byteenable                    (openmac_0_dma_byteenable),                   //                                      .byteenable
		.openmac_0_dma_read                          (openmac_0_dma_read),                         //                                      .read
		.openmac_0_dma_readdata                      (openmac_0_dma_readdata),                     //                                      .readdata
		.openmac_0_dma_readdatavalid                 (openmac_0_dma_readdatavalid),                //                                      .readdatavalid
		.openmac_0_dma_write                         (openmac_0_dma_write),                        //                                      .write
		.openmac_0_dma_writedata                     (openmac_0_dma_writedata),                    //                                      .writedata
		.pcp_0_cpu_bridge_address                    (pcp_0_cpu_bridge_address),                   //                      pcp_0_cpu_bridge.address
		.pcp_0_cpu_bridge_waitrequest                (pcp_0_cpu_bridge_waitrequest),               //                                      .waitrequest
		.pcp_0_cpu_bridge_burstcount                 (pcp_0_cpu_bridge_burstcount),                //                                      .burstcount
		.pcp_0_cpu_bridge_byteenable                 (pcp_0_cpu_bridge_byteenable),                //                                      .byteenable
		.pcp_0_cpu_bridge_read                       (pcp_0_cpu_bridge_read),                      //                                      .read
		.pcp_0_cpu_bridge_readdata                   (pcp_0_cpu_bridge_readdata),                  //                                      .readdata
		.pcp_0_cpu_bridge_readdatavalid              (pcp_0_cpu_bridge_readdatavalid),             //                                      .readdatavalid
		.pcp_0_cpu_bridge_write                      (pcp_0_cpu_bridge_write),                     //                                      .write
		.pcp_0_cpu_bridge_writedata                  (pcp_0_cpu_bridge_writedata),                 //                                      .writedata
		.pcp_0_cpu_bridge_debugaccess                (pcp_0_cpu_bridge_debugaccess),               //                                      .debugaccess
		.sram_0_uas_address                          (mm_interconnect_1_sram_0_uas_address),       //                            sram_0_uas.address
		.sram_0_uas_write                            (mm_interconnect_1_sram_0_uas_write),         //                                      .write
		.sram_0_uas_read                             (mm_interconnect_1_sram_0_uas_read),          //                                      .read
		.sram_0_uas_readdata                         (mm_interconnect_1_sram_0_uas_readdata),      //                                      .readdata
		.sram_0_uas_writedata                        (mm_interconnect_1_sram_0_uas_writedata),     //                                      .writedata
		.sram_0_uas_burstcount                       (mm_interconnect_1_sram_0_uas_burstcount),    //                                      .burstcount
		.sram_0_uas_byteenable                       (mm_interconnect_1_sram_0_uas_byteenable),    //                                      .byteenable
		.sram_0_uas_readdatavalid                    (mm_interconnect_1_sram_0_uas_readdatavalid), //                                      .readdatavalid
		.sram_0_uas_waitrequest                      (mm_interconnect_1_sram_0_uas_waitrequest),   //                                      .waitrequest
		.sram_0_uas_lock                             (mm_interconnect_1_sram_0_uas_lock),          //                                      .lock
		.sram_0_uas_debugaccess                      (mm_interconnect_1_sram_0_uas_debugaccess)    //                                      .debugaccess
	);

	soc_system_mm_interconnect_2 mm_interconnect_2 (
		.clk50_clk_clk                                                   (clk50_clk),                                                            //                                                 clk50_clk.clk
		.epcs_flash_controller_reset_reset_bridge_in_reset_reset         (rst_controller_006_reset_out_reset),                                   //         epcs_flash_controller_reset_reset_bridge_in_reset.reset
		.pcp_0_flash_bridge_translator_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                       // pcp_0_flash_bridge_translator_reset_reset_bridge_in_reset.reset
		.pcp_0_rst_clk50_reset_bridge_in_reset_reset                     (rst_controller_reset_out_reset),                                       //                     pcp_0_rst_clk50_reset_bridge_in_reset.reset
		.pcp_0_flash_bridge_address                                      (pcp_0_flash_bridge_address),                                           //                                        pcp_0_flash_bridge.address
		.pcp_0_flash_bridge_waitrequest                                  (pcp_0_flash_bridge_waitrequest),                                       //                                                          .waitrequest
		.pcp_0_flash_bridge_burstcount                                   (pcp_0_flash_bridge_burstcount),                                        //                                                          .burstcount
		.pcp_0_flash_bridge_byteenable                                   (pcp_0_flash_bridge_byteenable),                                        //                                                          .byteenable
		.pcp_0_flash_bridge_read                                         (pcp_0_flash_bridge_read),                                              //                                                          .read
		.pcp_0_flash_bridge_readdata                                     (pcp_0_flash_bridge_readdata),                                          //                                                          .readdata
		.pcp_0_flash_bridge_readdatavalid                                (pcp_0_flash_bridge_readdatavalid),                                     //                                                          .readdatavalid
		.pcp_0_flash_bridge_write                                        (pcp_0_flash_bridge_write),                                             //                                                          .write
		.pcp_0_flash_bridge_writedata                                    (pcp_0_flash_bridge_writedata),                                         //                                                          .writedata
		.pcp_0_flash_bridge_debugaccess                                  (pcp_0_flash_bridge_debugaccess),                                       //                                                          .debugaccess
		.epcs_flash_controller_epcs_control_port_address                 (mm_interconnect_2_epcs_flash_controller_epcs_control_port_address),    //                   epcs_flash_controller_epcs_control_port.address
		.epcs_flash_controller_epcs_control_port_write                   (mm_interconnect_2_epcs_flash_controller_epcs_control_port_write),      //                                                          .write
		.epcs_flash_controller_epcs_control_port_read                    (mm_interconnect_2_epcs_flash_controller_epcs_control_port_read),       //                                                          .read
		.epcs_flash_controller_epcs_control_port_readdata                (mm_interconnect_2_epcs_flash_controller_epcs_control_port_readdata),   //                                                          .readdata
		.epcs_flash_controller_epcs_control_port_writedata               (mm_interconnect_2_epcs_flash_controller_epcs_control_port_writedata),  //                                                          .writedata
		.epcs_flash_controller_epcs_control_port_chipselect              (mm_interconnect_2_epcs_flash_controller_epcs_control_port_chipselect)  //                                                          .chipselect
	);

	soc_system_irq_mapper irq_mapper (
		.clk           (clk50_clk),                      //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (pcp_0_sync_irq_irq)              //    sender.irq
	);

	soc_system_irq_mapper irq_mapper_001 (
		.clk           (clk50_clk),                      //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_001_receiver0_irq),   // receiver0.irq
		.sender_irq    (pcp_0_mac_irq_irq)               //    sender.irq
	);

	soc_system_irq_mapper_002 irq_mapper_002 (
		.clk           (clk50_clk),                      //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_002_receiver0_irq),   // receiver0.irq
		.sender_irq    (pcp_0_gp_irq_irq)                //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.reset_in1      (~reset_reset_n),                 // reset_in1.reset
		.reset_in2      (~reset_reset_n),                 // reset_in2.reset
		.clk            (clk50_clk),                      //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (~reset_reset_n),                     // reset_in1.reset
		.reset_in2      (~reset_reset_n),                     // reset_in2.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (~reset_reset_n),                     // reset_in1.reset
		.reset_in2      (~reset_reset_n),                     // reset_in2.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (~reset_reset_n),                     // reset_in1.reset
		.reset_in2      (~reset_reset_n),                     // reset_in2.reset
		.clk            (clk100_clk),                         //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (~reset_reset_n),                     // reset_in1.reset
		.reset_in2      (~reset_reset_n),                     // reset_in2.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_005 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (~reset_reset_n),                     // reset_in1.reset
		.reset_in2      (~reset_reset_n),                     // reset_in2.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_005_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (4),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_006 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (~reset_reset_n),                         // reset_in1.reset
		.reset_in2      (~reset_reset_n),                         // reset_in2.reset
		.reset_in3      (pcp_0_jtag_reset_reset),                 // reset_in3.reset
		.clk            (clk50_clk),                              //       clk.clk
		.reset_out      (rst_controller_006_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_006_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
